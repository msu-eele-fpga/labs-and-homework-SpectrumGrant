


entity synchronizer is
	port (
		clk	: in	std_ulogic;
		async	: in	std_ulogic;
		sync	: out	std_ulogic
	);
	
	
	